** sch_path: /home/thaonguyen06/eda/180mcuC/dls_nand_tran.sch
**.subckt dls_nand_tran
Vdd VDD GND 0.4
.save i(vdd)
Vin2 VinA GND pulse(0 0.4 0.5 0 0 5 10)
.save i(vin2)
Vin1 VinB GND pulse(0 0.4 0 0 0 5 10)
.save i(vin1)
X1 VinA VinB VDD GND Vout dls_nand
**** begin user architecture code


.include /home/thaonguyen06/eda/uniccass/share/pdk/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/thaonguyen06/eda/uniccass/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.tran 1s 50s
.save all

**** end user architecture code
**.ends

* expanding   symbol:  /home/thaonguyen06/eda/180mcuC/dls_nand.sym # of pins=5
** sym_path: /home/thaonguyen06/eda/180mcuC/dls_nand.sym
** sch_path: /home/thaonguyen06/eda/180mcuC/dls_nand.sch
.subckt dls_nand A B VP VN Y
*.iopin VP
*.ipin A
*.ipin B
*.iopin VN
*.opin Y
XM2 Y A net2 VP pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM1 Y A net1 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net1 B net3 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 Y B net2 VP pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 VN Y net3 VN pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 VP Y net2 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
